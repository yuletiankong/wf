`ifndef TEST_PARAMS_SVH
`define TEST_PARAMS_SVH

`define NUM_TESTS 300
`define NUM_TESTS_DEEP 200
`define INPUT_DIR "input_vectors"
`define OUTPUT_DIR "output"
`define SORTED_DIR "sorted_vectors"

`endif // TEST_PARAMS_SVH
